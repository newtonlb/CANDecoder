// Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
// Your use of Altera Corporation's design tools, logic functions 
// and other software and tools, and its AMPP partner logic 
// functions, and any output files from any of the foregoing 
// (including device programming or simulation files), and any 
// associated documentation or information are expressly subject 
// to the terms and conditions of the Altera Program License 
// Subscription Agreement, the Altera Quartus II License Agreement,
// the Altera MegaCore Function License Agreement, or other 
// applicable license agreement, including, without limitation, 
// that your use is for the sole purpose of programming logic 
// devices manufactured by Altera and sold by Altera or its 
// authorized distributors.  Please refer to the applicable 
// agreement for further details.

// Generated by Quartus II Version 15.0.0 Build 145 04/22/2015 SJ Web Edition
// Created on Wed Jun 14 03:48:00 2017

// synthesis message_off 10175

`timescale 1ns/1ps

module teste2 (input can_data, 
input sample,
output reg [10:0] bit_id_11 =11'bz,
output reg [28:0] bit_id_29 = 29'bz,
output reg [1:0] srr_rtr_ide = 0,
output reg data_frame = 0,
output reg getframe = 0,
output reg ext_frame = 0,
output reg std_frame = 0,
output reg rtr_ext = 1'bz,
output reg remote_frame = 0,
output reg [3:0] data_size
);

    /*input reset;
    input clock;
    input input1; //start of frame
    input input2;
    tri0 reset;
    tri0 input1;
    tri0 input2;
    reg [2:0] fstate; // estado atual
	reg [7:0] state=0;
    reg [2:0] reg_fstate; // próximo estado
    parameter state1=0,state2=1,state3=2;
	*/ 
	reg [28:0] arbitration_field = 0; 
	
	reg[7:0] state = 0;
	reg [9:0] count = 0; //vai contar os bits do Arbitration Field
	reg s0;
	reg r0;
	reg r1;
	reg r2;
	
    

    always @(posedge sample)
    begin
        case (state)
                0 : begin
                    	if ((can_data == 0)) // start of frame
			begin
				state = 1;
				count = 29;
			
                    	
                    	
			end
			else //bit 1
			begin
				state = 0;
				count = count + 1;
				if(count == 6)
				begin
					$display ("deu erro");//vai dar erro aqui pq veio 6 bits 1
				end
			end
				
                        
                end
                1 : begin
			state = 1;
			arbitration_field[count-1] = can_data;
			count = count -1;
			if(count == 18) // pegou os 11 bits
			begin
				state = 2;
				count = 2;
			end
                    	 // Acabou o Arbitration Field
                        
                    	// Inserting 'else' block to prevent latch inference
                end
                2 : begin
                    	srr_rtr_ide[count -1] = can_data;
			count = count -1;
			if(count == 0)
			begin
				if(srr_rtr_ide == 2'b00)// � um frame de dados, 11 bits
				
				begin
					$display ("� um frame de dados, 11 bits");
					bit_id_11 = arbitration_field[28:18];
					data_frame = 1;
					std_frame = 1;
					state = 5;

				end
				if(srr_rtr_ide == 2'b10)// � um frame remote request, 11 bits
				begin
					$display ("eh um remote request, 11 bits");
					bit_id_11 = arbitration_field[28:18];
					std_frame = 1;
					remote_frame = 1;
					state = 5;
					
				end
				if(srr_rtr_ide == 2'b11) //� o srr e � um frame de 29 bits
					
				begin
					$display ("eh um frame de 29 bits");
					bit_id_11 = arbitration_field[28:18];
					ext_frame = 1;
					count = 18;
					state = 3;
				
				end
               	 	end
		end
		
		3: begin //se for 29 bits, tem que pegar o resto do ID
		
		
			
			arbitration_field[count-1] = can_data;	
			count = count -1;
			
			if (count == 0) //terminou os 29-bits
			begin 
				bit_id_29[28:0] = arbitration_field[28:0];
				state = 4; //vai pegar o RTR do estendido
			end
			
				
				
		end

		4: begin //um estado s� pra pegar o rtr do estendido
			rtr_ext = can_data;
			if(rtr_ext == 0)
			begin
			$display("ele ta acusando que eh um data frame");
				data_frame = 1;
	      			//� um frame de dados estendido
			end
			if(rtr_ext == 1)
			begin
				remote_frame = 1;
				//� um remote frame estendido
			end
			state = 6; //pegar os dois bits reservados
			count = 2;

		
		end
		

		5: begin //tratar bit reservado frame dados
			r0 = can_data;
			count = 4;			
			state = 7;
		end
		
		6: begin //pegando os dois bits reservados do esetendido
			count = count -1;
			$display("can_data %h count %d", can_data, count);
			if (count == 0)
			begin
				state = 7;
				count = 4;
			end
			else
			begin
				state = 6;
			end

		end
		7: begin //pegar os 4 bits indicando a quantidade de bytes de dados
			data_size[count-1] = can_data;
			count = count -1;
			if(count == 0)
			begin
				//vai pegar os dados agora
				state = 8;
			end
		end

                8: begin
			getframe = 1;
		end
		default: begin
                    $display ("Reach undefined state");
                end
      endcase
    end
endmodule // teste2
